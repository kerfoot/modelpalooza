netcdf modelGliderFlatNc {
dimensions:
	time = 262 ;
	traj_strlen = 18 ;
variables:
	double time(time) ;
		time:ancillary_variables = " " ;
		time:long_name = "Time" ;
		time:standard_name = "time" ;
		time:units = "seconds since 1970-01-01T00:00:00Z" ;
	char trajectory(traj_strlen) ;
		trajectory:cf_role = "trajectory_id" ;
		trajectory:comment = "A trajectory is a glider deployment" ;
		trajectory:long_name = "Trajectory Name" ;
	double lat(time) ;
		lat:long_name = "Latitude" ;
		lat:standard_name = "latitude" ;
		lat:units = "degrees_north" ;
		lat:_FillValue = -999. ;
	double lon(time) ;
		lon:long_name = "Longitude" ;
		lon:standard_name = "longitude" ;
		lon:units = "degrees_east" ;
		lon:_FillValue = -999. ;
	double depth(time) ;
		depth:comment = " " ;
		depth:instrument = "instrument_ctd" ;
		depth:long_name = "Depth" ;
		depth:observation_type = "calculated" ;
		depth:positive = "down" ;
		depth:standard_name = "depth" ;
		depth:units = "meters" ;
		depth:valid_max = 2000. ;
		depth:valid_min = 0. ;
		depth:_FillValue = -999. ;
	double temperature(time) ;
		temperature:instrument = "instrument_ctd" ;
		temperature:long_name = "Temperature" ;
		temperature:observation_type = "measured" ;
		temperature:standard_name = "sea_water_temperature" ;
		temperature:units = "Celsius" ;
		temperature:valid_max = 40. ;
		temperature:valid_min = -5. ;
		temperature:_FillValue = -999. ;
	double salinity(time) ;
		salinity:instrument = "instrument_ctd" ;
		salinity:long_name = "Salinity" ;
		salinity:observation_type = "calculated" ;
		salinity:standard_name = "sea_water_practical_salinity" ;
		salinity:units = "1e-3" ;
		salinity:valid_max = 40. ;
		salinity:valid_min = 0. ;
		salinity:_FillValue = -999. ;
	double density(time) ;
		density:instrument = "instrument_ctd" ;
		density:long_name = "Density" ;
		density:observation_type = "calculated" ;
		density:standard_name = "sea_water_density" ;
		density:units = "kg m-3" ;
		density:valid_max = 1040. ;
		density:valid_min = 1015. ;
		density:_FillValue = -999. ;
    double u(time) ;
		u:long_name = "Eastward Sea Water Velocity" ;
		u:standard_name = "eastward_sea_water_velocity" ;
		u:units = "m s-1" ;
		u:_FillValue = -999. ;
    double v(time) ;
		v:long_name = "Northward Sea Water Velocity" ;
		v:standard_name = "northward_sea_water_velocity" ;
		v:units = "m s-1" ;
		v:_FillValue = -999. ;
	int profile_id ;
		profile_id:long_name = "Sequential Profile ID" ;
		profile_id:_FillValue = -127b ;
	double profile_time ;
		profile_time:long_name = "Profile Center Time" ;
		profile_time:standard_name = "time" ;
		profile_time:units = "seconds since 1970-01-01T00:00:00Z" ;
		profile_time:_FillValue = -999. ;
	double profile_lat ;
		profile_lat:long_name = "Profile Center Latitude" ;
		profile_lat:standard_name = "latitude" ;
		profile_lat:units = "degrees_north" ;
		profile_lat:_FillValue = -999. ;
	double profile_lon ;
		profile_lon:long_name = "Profile Center Longitude" ;
		profile_lon:standard_name = "longitude" ;
		profile_lon:units = "degrees_east" ;
		profile_lon:_FillValue = -999. ;

// global attributes:
		:Metadata_Conventions = "CF-1.6, Unidata Dataset Discovery v1.0" ;
		:Conventions = "CF-1.6" ;
		:acknowledgment = "Modeled profile data provided by the National Weather Service's National Centers for Environmental Prediction (NCEP).  Glider profile locations provided by the Rutgers University Coastal Ocean Observation Lab." ;
		:comment = " " ;
		:contributor_name = "John Kerfoot" ;
		:contributor_role = "Data Manager" ;
		:creator_email = "kerfoot@marine.rutgers.edu" ;
		:creator_name = "John Kerfoot" ;
		:creator_url = "http://marine.rutgers.edu/cool/auvs" ;
        :date_created = " " ;
        :date_issued = " " ;
		:date_modified = " " ;
		:format_version = "rtofsGliderFlatNc" ;
        :history = " " ;
		:id = " " ;
		:institution = "NCEP" ;
		:keywords = "Models, Government Agencies-U.S. Federal Agencies > DOC/NOAA/NWS/NCEP, National Centers for Environmental Prediction, National Weather Service, http://www.ncep.noaa.gov/, Oceans > Ocean Pressure > Water Pressure, Oceans > Ocean Temperature > Water Temperature, Oceans > Salinity/Density > Conductivity, Oceans > Salinity/Density > Density, Oceans > Salinity/Density > Salinity" ;
		:keywords_vocabulary = "GCMD Science Keywords" ;
		:license = "Rutgers University and NCEP assume no liability resulting from the use of these data. No data quality assurance steps have been implemented on this data to date.  These files are to be used for comparison with measured Slocum glider vertical profiles.  This dataset is represents a 'virtual' glider dataset sampled from RTOFS at each glider profile location." ;
		:metadata_link = " " ;
		:naming_authority = "edu.rutgers.marine" ;
		:platform_type = "Model" ;
        :processing_level = " " ;
		:project = "Modelpalooza" ;
		:publisher_email = "kerfoot@marine.rutgers.edu" ;
		:publisher_name = "John Kerfoot" ;
		:publisher_url = "http://marine.rutgers.edu/cool/auvs" ;
		:references = " " ;
		:sea_name = "South Atlantic Ocean" ;
		:source = "Global RTOFS model forecast" ;
		:standard_name_vocabulary = "CF-1.6" ;
		:summary = "The Global RTOFS ocean model is based on an eddy resolving 1/12 degree global HYCOM (HYbrid Coordinates Ocean Model) (Chassignet et al., 2009) and is part of a larger national backbone capability of ocean modeling at NWS in a strong partnership with US Navy. The Global RTOFS ocean model became operational 25 October 2011.  RTOFS vertical profiles are selected for the closest grid point to the measured glider GPS profile position. This dataset represents a 'virtual' glider dataset containing the closest modeled vertical profiles along the glider's path." ;
		:title = " " ;
}
